//7 to 128 bit decoder module
module decoder_7_128(input_7, output_128);
input [6:0] input_7;

output [127:0] output_128;

assign output_128 = (input_7 == 0) ? 128'h00000000000000000000000000000001 :
				(input_7 == 1) ? 128'h00000000000000000000000000000002 :
				(input_7 == 2) ? 128'h00000000000000000000000000000004 :
				(input_7 == 3) ? 128'h00000000000000000000000000000008 :
				(input_7 == 4) ? 128'h00000000000000000000000000000010 :
				(input_7 == 5) ? 128'h00000000000000000000000000000020 :
				(input_7 == 6) ? 128'h00000000000000000000000000000040 :
				(input_7 == 7) ? 128'h00000000000000000000000000000080 :
				(input_7 == 8) ? 128'h00000000000000000000000000000100 :
				(input_7 == 9) ? 128'h00000000000000000000000000000200 :
				(input_7 == 10) ? 128'h00000000000000000000000000000400 :
				(input_7 == 11) ? 128'h00000000000000000000000000000800 :
				(input_7 == 12) ? 128'h00000000000000000000000000001000 :
				(input_7 == 13) ? 128'h00000000000000000000000000002000 :
				(input_7 == 14) ? 128'h00000000000000000000000000004000 :
				(input_7 == 15) ? 128'h00000000000000000000000000008000 :
				(input_7 == 16) ? 128'h00000000000000000000000000010000 :
				(input_7 == 17) ? 128'h00000000000000000000000000020000 :
				(input_7 == 18) ? 128'h00000000000000000000000000040000 :
				(input_7 == 19) ? 128'h00000000000000000000000000080000 :
				(input_7 == 20) ? 128'h00000000000000000000000000100000 :
				(input_7 == 21) ? 128'h00000000000000000000000000200000 :
				(input_7 == 22) ? 128'h00000000000000000000000000400000 :
				(input_7 == 23) ? 128'h00000000000000000000000000800000 :
				(input_7 == 24) ? 128'h00000000000000000000000001000000 :
				(input_7 == 25) ? 128'h00000000000000000000000002000000 :
				(input_7 == 26) ? 128'h00000000000000000000000004000000 :
				(input_7 == 27) ? 128'h00000000000000000000000008000000 :
				(input_7 == 28) ? 128'h00000000000000000000000010000000 :
				(input_7 == 29) ? 128'h00000000000000000000000020000000 :
				(input_7 == 30) ? 128'h00000000000000000000000040000000 :
				(input_7 == 31) ? 128'h00000000000000000000000080000000 :
				(input_7 == 32) ? 128'h00000000000000000000000100000000 :
				(input_7 == 33) ? 128'h00000000000000000000000200000000 :
				(input_7 == 34) ? 128'h00000000000000000000000400000000 :
				(input_7 == 35) ? 128'h00000000000000000000000800000000 :
				(input_7 == 36) ? 128'h00000000000000000000001000000000 :
				(input_7 == 37) ? 128'h00000000000000000000002000000000 :
				(input_7 == 38) ? 128'h00000000000000000000004000000000 :
				(input_7 == 39) ? 128'h00000000000000000000008000000000 :
				(input_7 == 40) ? 128'h00000000000000000000010000000000 :
				(input_7 == 41) ? 128'h00000000000000000000020000000000 :
				(input_7 == 42) ? 128'h00000000000000000000040000000000 :
				(input_7 == 43) ? 128'h00000000000000000000080000000000 :
				(input_7 == 44) ? 128'h00000000000000000000100000000000 :
				(input_7 == 45) ? 128'h00000000000000000000200000000000 :
				(input_7 == 46) ? 128'h00000000000000000000400000000000 :
				(input_7 == 47) ? 128'h00000000000000000000800000000000 :
				(input_7 == 48) ? 128'h00000000000000000001000000000000 :
				(input_7 == 49) ? 128'h00000000000000000002000000000000 :
				(input_7 == 50) ? 128'h00000000000000000004000000000000 :
				(input_7 == 51) ? 128'h00000000000000000008000000000000 :
				(input_7 == 52) ? 128'h00000000000000000010000000000000 :
				(input_7 == 53) ? 128'h00000000000000000020000000000000 :
				(input_7 == 54) ? 128'h00000000000000000040000000000000 :
				(input_7 == 55) ? 128'h00000000000000000080000000000000 :
				(input_7 == 56) ? 128'h00000000000000000100000000000000 :
				(input_7 == 57) ? 128'h00000000000000000200000000000000 :
				(input_7 == 58) ? 128'h00000000000000000400000000000000 :
				(input_7 == 59) ? 128'h00000000000000000800000000000000 :
				(input_7 == 60) ? 128'h00000000000000001000000000000000 :
				(input_7 == 61) ? 128'h00000000000000002000000000000000 :
				(input_7 == 62) ? 128'h00000000000000004000000000000000 :
				(input_7 == 63) ? 128'h00000000000000008000000000000000 :
				(input_7 == 64) ? 128'h00000000000000010000000000000000 :
				(input_7 == 65) ? 128'h00000000000000020000000000000000 :
				(input_7 == 66) ? 128'h00000000000000040000000000000000 :
				(input_7 == 67) ? 128'h00000000000000080000000000000000 :
				(input_7 == 68) ? 128'h00000000000000100000000000000000 :
				(input_7 == 69) ? 128'h00000000000000200000000000000000 :
				(input_7 == 70) ? 128'h00000000000000400000000000000000 :
				(input_7 == 71) ? 128'h00000000000000800000000000000000 :
				(input_7 == 72) ? 128'h00000000000001000000000000000000 :
				(input_7 == 73) ? 128'h00000000000002000000000000000000 :
				(input_7 == 74) ? 128'h00000000000004000000000000000000 :
				(input_7 == 75) ? 128'h00000000000008000000000000000000 :
				(input_7 == 76) ? 128'h00000000000010000000000000000000 :
				(input_7 == 77) ? 128'h00000000000020000000000000000000 :
				(input_7 == 78) ? 128'h00000000000040000000000000000000 :
				(input_7 == 79) ? 128'h00000000000080000000000000000000 :
				(input_7 == 80) ? 128'h00000000000100000000000000000000 :
				(input_7 == 81) ? 128'h00000000000200000000000000000000 :
				(input_7 == 82) ? 128'h00000000000400000000000000000000 :
				(input_7 == 83) ? 128'h00000000000800000000000000000000 :
				(input_7 == 84) ? 128'h00000000001000000000000000000000 :
				(input_7 == 85) ? 128'h00000000002000000000000000000000 :
				(input_7 == 86) ? 128'h00000000004000000000000000000000 :
				(input_7 == 87) ? 128'h00000000008000000000000000000000 :
				(input_7 == 88) ? 128'h00000000010000000000000000000000 :
				(input_7 == 89) ? 128'h00000000020000000000000000000000 :
				(input_7 == 90) ? 128'h00000000040000000000000000000000 :
				(input_7 == 91) ? 128'h00000000080000000000000000000000 :
				(input_7 == 92) ? 128'h00000000100000000000000000000000 :
				(input_7 == 93) ? 128'h00000000200000000000000000000000 :
				(input_7 == 94) ? 128'h00000000400000000000000000000000 :
				(input_7 == 95) ? 128'h00000000800000000000000000000000 :
				(input_7 == 96) ? 128'h00000001000000000000000000000000 :
				(input_7 == 97) ? 128'h00000002000000000000000000000000 :
				(input_7 == 98) ? 128'h00000004000000000000000000000000 :
				(input_7 == 99) ? 128'h00000008000000000000000000000000 :
				(input_7 == 100) ? 128'h00000010000000000000000000000000 :
				(input_7 == 101) ? 128'h00000020000000000000000000000000 :
				(input_7 == 102) ? 128'h00000040000000000000000000000000 :
				(input_7 == 103) ? 128'h00000080000000000000000000000000 :
				(input_7 == 104) ? 128'h00000100000000000000000000000000 :
				(input_7 == 105) ? 128'h00000200000000000000000000000000 :
				(input_7 == 106) ? 128'h00000400000000000000000000000000 :
				(input_7 == 107) ? 128'h00000800000000000000000000000000 :
				(input_7 == 108) ? 128'h00001000000000000000000000000000 :
				(input_7 == 109) ? 128'h00002000000000000000000000000000 :
				(input_7 == 110) ? 128'h00004000000000000000000000000000 :
				(input_7 == 111) ? 128'h00008000000000000000000000000000 :
				(input_7 == 112) ? 128'h00010000000000000000000000000000 :
				(input_7 == 113) ? 128'h00020000000000000000000000000000 :
				(input_7 == 114) ? 128'h00040000000000000000000000000000 :
				(input_7 == 115) ? 128'h00080000000000000000000000000000 :
				(input_7 == 116) ? 128'h00100000000000000000000000000000 :
				(input_7 == 117) ? 128'h00200000000000000000000000000000 :
				(input_7 == 118) ? 128'h00400000000000000000000000000000 :
				(input_7 == 119) ? 128'h00800000000000000000000000000000 :
				(input_7 == 120) ? 128'h01000000000000000000000000000000 :
				(input_7 == 121) ? 128'h02000000000000000000000000000000 :
				(input_7 == 122) ? 128'h04000000000000000000000000000000 :
				(input_7 == 123) ? 128'h08000000000000000000000000000000 :
				(input_7 == 124) ? 128'h10000000000000000000000000000000 :
				(input_7 == 125) ? 128'h20000000000000000000000000000000 :
				(input_7 == 126) ? 128'h40000000000000000000000000000000 :
				(input_7 == 127) ? 128'h80000000000000000000000000000000 :
				128'hxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
endmodule
